module stage_mem(
);

endmodule
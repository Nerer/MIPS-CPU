module register();